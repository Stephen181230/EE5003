module tb();

// 16 bits potential width 
// 16 bits weight width 
// 16 bits range(-32768,32767)
// width memory depth = 32
// 
parameter I_I = 8; //reg width for I
parameter I_J = 8; //reg width for J
parameter I_K = 8; //reg width for K
parameter I_T = 8; //reg width for L
parameter K_I             = 8; //reg width for kernel I
parameter K_J             = 8; //reg width for kernel J
parameter K_K             = 1;
parameter MAX_KERNEL_NUM  = 16;//max kernel num
parameter BASE_ADDR_WIDTH = 32;
parameter DEPTH           = 16; // for input fifo DEPTH
parameter WIDTH           = 32; // for input fifo WIDTH
parameter i_width         = 8;
parameter j_width         = 8;
parameter k_width         = 8;
parameter l_width         = 8;
parameter WEIGHT_WIDTH    = 32;// 16 signed reg
parameter POTENTIAL_WIDTH = 32;// poential memory width
parameter WEIGHT_DEPTH    = 32; 
parameter POTENTIAL_DEPTH = 16;
parameter NUM_ARB         = 6;
parameter PE_NUM          = 4;
parameter POST_WIDTH      = 32;


  //Ports
  reg  potential_read_en; 
  reg  potential_write_en; 
  reg [$clog2(POTENTIAL_DEPTH)-1:0] potential_raddr_cluster; //addr no need to signed reg
  reg [$clog2(POTENTIAL_DEPTH)-1:0] potential_waddr_cluster; //addr no need to signed reg
  reg signed [POTENTIAL_WIDTH*MAX_KERNEL_NUM-1:0] potential_wdata_cluster; // write data need signed reg
  reg  clk;
  reg  rst;
  reg [PE_NUM-1:0] start;
  reg start_sche;
  reg signed [POTENTIAL_WIDTH-1:0] threhold;
  reg signed [POTENTIAL_WIDTH-1:0] rest_value;
  reg [2:0]working_mode;
  reg [31:0] w_data;
  reg [31:0] w_value;
  reg [PE_NUM-1:0] w_mem_wen;
  reg [WEIGHT_WIDTH*MAX_KERNEL_NUM-1:0] w_mem_wdata;
  reg [$clog2(WEIGHT_DEPTH)-1:0] w_mem_waddr;
  reg [K_I-1:0] k_i;
  reg [K_J-1:0] k_j;
  reg [I_I-1:0] i_i;
  reg [I_J-1:0] i_j;
  reg [BASE_ADDR_WIDTH-1:0] base_addr;
  reg pre_grant;
  reg post_grant;
  reg signed [WEIGHT_WIDTH-1:0]weight_inst;
  reg [POST_WIDTH-1:0] post_addr;
  reg [15:0]output_neuron_num;
  reg [I_T-1:0] timestamp;
  wire [POST_WIDTH-1:0] post_waddr;
  wire signed [POST_WIDTH-1:0] post_wdata;
  wire [PE_NUM-1:0] finish;
  wire [NUM_ARB-1:0] Read_req;
  wire [NUM_ARB-1:0] Write_req;
  wire [NUM_ARB-1:0] Read_grant;
  wire  post_req;
  wire [3:0] PE_grant;
  wire [4*$clog2(POTENTIAL_DEPTH)-1:0]  potential_raddr;
  wire [4*$clog2(POTENTIAL_DEPTH)-1:0]  potential_waddr;
  wire flagout;
  wire [$clog2(DEPTH)-1:0]          Write_Addr;
  wire [$clog2(DEPTH)-1:0]          Read_Addr;
  wire signed[POTENTIAL_WIDTH*MAX_KERNEL_NUM-1:0]      Read_data;
  wire finish_sche;


  



  cluster # (
    .I_I(I_I),
    .I_J(I_J),
    .I_K(I_K),
    .K_I(K_I),
    .K_J(K_J),
    .K_K(K_K),
    .BASE_ADDR_WIDTH(BASE_ADDR_WIDTH),
    .DEPTH(DEPTH),
    .WIDTH(WIDTH),
    .i_width(i_width),
    .j_width(j_width),
    .k_width(k_width),
    .l_width(l_width),
    .WEIGHT_WIDTH(WEIGHT_WIDTH),
    .POTENTIAL_WIDTH(POTENTIAL_WIDTH),
    .WEIGHT_DEPTH(WEIGHT_DEPTH),
    .POTENTIAL_DEPTH(POTENTIAL_DEPTH),
    .NUM_ARB(NUM_ARB),
    .PE_NUM(PE_NUM),
    .POST_WIDTH(POST_WIDTH),
    .MAX_KERNEL_NUM(MAX_KERNEL_NUM)
  )
  cluster_inst (
    .potential_read_en(potential_read_en),
    .potential_write_en(potential_write_en),
    .potential_raddr_cluster(potential_raddr_cluster),
    .potential_waddr_cluster(potential_waddr_cluster),
    .potential_wdata_cluster(potential_wdata_cluster),
    .clk(clk),
    .rst(rst),
    .start(start),
    .threhold(threhold),
    .rest_value(rest_value),
    .working_mode(working_mode),
    .w_data(w_data),
    .w_mem_wen(w_mem_wen),
    .w_mem_wdata(w_mem_wdata),
    .w_mem_waddr(w_mem_waddr),
    .k_i(k_i),
    .k_j(k_j),
    .i_i(i_i),
    .i_j(i_j),
    .base_addr(base_addr),
    .pre_grant(pre_grant),
    .post_grant(post_grant),
    .post_addr(post_addr),
    .post_waddr(post_waddr),
    .post_wdata(post_wdata),
    .finish(finish),
    .post_req(post_req),
    .Potential_raddr(potential_raddr),
    .Potential_waddr(potential_waddr),
    .Read_req(Read_req),
    .Write_req(Write_req),
    .Read_grant(Read_grant),
    .flagout(flagout),
    .Write_Addr       (Write_Addr),
    .Read_Addr        (Read_Addr),
    .PE_grant         (PE_grant),
    .Read_data         (Read_data),
    .output_neuron_num (output_neuron_num),
    .finish_sche      (finish_sche),
    .timestamp        (timestamp),
    .w_value          (w_value),
    .start_sche       (start_sche)

    
  );

  initial begin
    potential_read_en = 0;
    potential_write_en = 0; 
    potential_raddr_cluster = 0;
    potential_waddr_cluster = 0;
    potential_wdata_cluster = 0;
    clk  = 0;
    rst             =0;
    start           =0;
    threhold        =32'b0000_0000_0000_0000_1000_0000_0000_0000;
    rest_value      =0;
    working_mode    =3'b010;
    w_data          =0;
    w_mem_wen       =0;      
    w_mem_wdata     =0;  
    w_mem_waddr     =0;
    k_i             =0;
    k_j             =0;
    i_i             =0;
    i_j             =0;
    base_addr       =0;
    post_grant      =1;
    pre_grant           =0;
    post_addr       =0;
    output_neuron_num = 10;
    weight_inst     =0;
    timestamp       =0;
    start_sche      =0;

    

    #20 //write weight PE=1
    rst =1;
    k_i =0;
    k_j =0;
    i_i =0;
    i_j =0;
    w_mem_wen = 4'b0001;
    w_mem_waddr      =0; //neuron ID = 0
    w_mem_wdata = 512'b00000000000000001101111010010010000000000000000000001101101111010000000000000000011101011000101011111111111111110000100000011011000000000000000000010100110100010000000000000000001000110011010000000000000000001111111010110010000000000000000011010110011100011111111111111111001111101000111111111111111111110101100100001101000000000000000011110111101101101111111111111111011001001001000000000000000000001110001000100001111111111111111100000101100101011111111111111111010001010111100011111111111111110111101110010000;
    #20
    w_mem_waddr = 1; //neuron ID = 4
    w_mem_wdata = 512'b00000000000000001010010101010110000000000000000001001101101111100000000000000000101011101011101111111111111111110111110111100011111111111111111100001011100111010000000000000000100001010101111011111111111111110000111111000110111111111111111111100001110111110000000000000000101101000000110000000000000000001011100111101100000000000000000001000011111101001111111111111111101100100101110100000000000000001110111101111001111111111111111101011110001101111111111111111111000111000000001111111111111111110001111000010000;
    
    #20
    w_mem_waddr = 2; //neuron ID = 8
    w_mem_wdata = 512'b00000000000000000100010101010111000000000000000001010111100010011111111111111111110100111101011100000000000000000000001100001001000000000000000000010000011011110000000000000000110101001000011111111111111111111001011010011101000000000000000011100100100110010000000000000000100101001101001011111111111111111000111010110010000000000000000010011010111011010000000000000000100101111001111111111111111111111111101100010100111111111111111100000100010011101111111111111111000101011111001111111111111111110000101110010001;


    
    #20 //write weight PE=1
    w_mem_wen = 4'b0010;
    w_mem_waddr      =0; //neuron ID = 1
    w_mem_wdata = 512'b00000000000000000101010010010110111111111111111101010001110010011111111111111111110100111010001111111111111111111011010111101011111111111111111110001101101001001111111111111111110000000010101100000000000000000111110101100100000000000000000001111101011010101111111111111111100100111110001011111111111111111111001001110011000000000000000001111100111001000000000000000000101111100000010011111111111111111001001101100101111111111111111111011100110110001111111111111111000000111010011000000000000000001011001110010100;
    
    #20
    w_mem_waddr      =1; //neuron ID = 5
    w_mem_wdata = 512'b11111111111111110010000010001010111111111111111111001111000000010000000000000000010001001101111111111111111111110111110101100001111111111111111100001100101110101111111111111111001011100001000000000000000000001101011101110111111111111111111101111000001111111111111111111111001001000110101011111111111111111110111100100111111111111111111101000001010100010000000000000000111000111110001000000000000000000011101100111001000000000000000010100010110011111111111111111111111110110101001011111111111111110011011110000000;
    #20
    w_mem_waddr = 2; //neuron ID = 9
    w_mem_wdata = 512'b00000000000000001010011100100100000000000000000011101110100001000000000000000000110011001000101100000000000000001100000001100001000000000000000010001000010000111111111111111111010011001101111100000000000000000011110101010001111111111111111100110010111110111111111111111111100001000010110100000000000000001100100100000110000000000000000001101110001111000000000000000000000100001000010011111111111111111010101100011010111111111111111110010101101101011111111111111111000110101001110000000000000000001010110001110111;
        
    #20 //write weight PE=1
    w_mem_wen = 4'b0100;
    w_mem_waddr      =0; //neuron ID = 2
    w_mem_wdata = 512'b00000000000000001111110010100110111111111111111101010000000000101111111111111111011000001010100111111111111111111110010111110110000000000000000010110000001100101111111111111111011010111100110111111111111111110111000001000111111111111111111110111110111011101111111111111111001000001010011011111111111111110111111111011101111111111111111100011001001111010000000000000000101000100000010100000000000000001100011110110100111111111111111110001001100000010000000000000000100111000101010011111111111111111001011000011010;
    
    #20
    w_mem_waddr      =1; //neuron ID = 6
    w_mem_wdata = 512'b11111111111111110101001001110100000000000000000000000010110111011111111111111111100100000111001100000000000000000110000010110110000000000000000000110000011001100000000000000000111000100100111011111111111111111001000000001010000000000000000010110010000111001111111111111111000011000011010011111111111111110100100000000110111111111111111110110111010000110000000000000000001111100111001000000000000000000000101001001011000000000000000011010010001110111111111111111111001000101100111111111111111111110100101100110011;
    
    #20 //write weight PE=1
    rst =1;
    w_mem_wen = 4'b1000;
    w_mem_waddr      =0; //neuron ID = 3
    w_mem_wdata = 512'b00000000000000000011111010111001111111111111111101110100111110101111111111111111001000101100111111111111111111111010101110010110000000000000000010101100001111001111111111111111101110101000101100000000000000000011110010001011000000000000000001000010011010001111111111111111111100011110010000000000000000001110100100101011111111111111111111001100011010000000000000000000100001010011000011111111111111111010010010101101000000000000000010111000100101110000000000000000010001111000000000000000000000000111101010001100;    
    
    #20
    w_mem_waddr      =1; //neuron ID = 7
    w_mem_wdata = 512'b00000000000000000001001001100111000000000000000000111010100000101111111111111111100110110010001100000000000000001000001001110001000000000000000001011101000011011111111111111111000100111010000000000000000000000010111011111111000000000000000001011100100010110000000000000000110011111001110111111111111111110000100100000111000000000000000010001110010100011111111111111111111101011010001000000000000000001100000000010110111111111111111101000001000101110000000000000000000001011111010000000000000000001111110101011010;    
    

    

    #20 //write input 
    w_mem_wen       =0;
    w_mem_waddr     =0;
    w_mem_wdata     =0;
    
    #20
    start = 4'b1111;
    pre_grant      =1;
    w_data          =0; //neuron id = 0
    w_value         =2;

    
    #60 //write input 
    w_data          =1; //neuron id = 1
    w_value         =2;
//    #20
//    w_data          =32'b00_00000_00000_00010_00001_00010_00000; //i=1, j=0, k=2
    
    #60 //write input 
    w_data          =2;
    w_value         =2;
    
    #60 //write input 
    w_data          =3;
    w_value         =2;
    
//    #60 //write input 
//    w_data          =9;


    #60
    w_data =0;
    pre_grant =0;
    

    #500
    start_sche = 1;

    
    

    

    

    
    


    
  end
always #10  clk = ! clk ;

endmodule

